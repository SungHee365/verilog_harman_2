`timescale 1ns / 1ps

module rom (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:32];

    initial begin
        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ opcode; // L-Type
        rom[0] = 32'b000000000100_00000_000_00011_0000011; // lb x2, 4(x0); [0:7]
        rom[1] = 32'b000000000100_00000_001_00011_0000011; // lh x3, 4(x0); [0:15]
        rom[2] = 32'b000000000100_00000_010_00011_0000011; // lw x4, 4(x0); [0:31]
        rom[3] = 32'b000000000100_00000_100_00011_0000011; // lbu x5, 4(x0); [0:7] // rdata 분할해야됨 5가지 종류로
        rom[4] = 32'b000000000100_00000_101_00011_0000011; // lhu x6, 4(x0); [0:15]
    end
    assign data = rom[addr[31:2]];
endmodule

/*
    initial begin
        
        //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _opcode; // R-Type
        rom[0] = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x2, x1      
        rom[1] = 32'b0100000_00001_00010_000_00101_0110011; // sub x5, x2, x1
        //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ opcode; // S-Type
        rom[2] = 32'b0000000_00010_00000_010_01000_0100011; // sw x2, 8(x0);
        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ opcode; // L-Type
        rom[3] = 32'b000000001000_00000_010_00011_0000011; // lw x3, 8(x0);
        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ opcode; // I-Type
        rom[4] = 32'b000000001000_00010_000_00110_0010011; // addi x6, x2, 8
        //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ opcode // B-Type
        rom[5] = 32'b0000000_00001_00001_000_11100_1100011;

        //테스트용
        //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _opcode; // R-Type
        rom[0] = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x2, x1 12+11=23      
        rom[1] = 32'b0100000_00001_00010_000_00101_0110011; // sub x5, x2, x1 12-11=1
        rom[2] = 32'b0000000_00101_00101_001_00110_0110011; // sll x6, x5, x5 1 << 1   = 2
        rom[3] = 32'b0000000_00101_00101_101_00111_0110011; // srl x7, x5, x5 1 >> 1   = 0
        rom[4] = 32'b0100000_00011_00001_000_01000_0110011; // sub x8, x1, x3 11 - 13  = -2
        rom[5] = 32'b0100000_00110_01000_101_01001_0110011; // sra x9, x8, x5 -2 >>> 1 = -1
        rom[6] = 32'b0000000_01000_00110_010_01010_0110011; // slt x10,x6, x8  2 < -2  = 0
        rom[7] = 32'b0000000_01000_00110_011_01011_0110011; // sltu x11,x6, x8         = 1
        rom[8] = 32'b0000000_00110_00101_100_01100_0110011; // xor x12,x5, x6 2 ^ 1    = 3
        rom[9] = 32'b0000000_00111_00101_110_01101_0110011; // or  x13,x5, x7 1 | 0    = 1
        rom[10] = 32'b0000000_00111_00101_111_01110_0110011; //and x14,x5, x7 1 & 0    = 0
        //rom[x]= 32'b imm12      _ rs1 _f3 _ rd  _ opcode; // I-Type
        rom[11] = 32'b000000000100_00111_000_01111_0010011; //addi x15, x7, 0 + 4 = 4
        rom[12] = 32'b111111111110_00111_010_10000_0010011; //slti x16, x7, 0 < -2 = 0
        rom[13] = 32'b111111111110_00111_011_10001_0010011; //sltiu x17, x7, 0 < ?? = 1
        rom[14] = 32'b000000000001_00110_100_10010_0010011; //xori x18, x6, 2 ^ 1 = 3
        rom[15] = 32'b000000000001_00110_110_10011_0010011; // ori x19, x6, 2 | 1 = 3
        rom[16] = 32'b000000000001_00110_111_10100_0010011; // and x20, x6, 2 & 1 = 0 
        rom[17] = 32'b000000000001_00110_001_10101_0010011; // slli x21, x6, 2 << 1 = 4
        rom[18] = 32'b000000000001_00110_101_10110_0010011; // srli x22, x6  2 >> 1 = 1
        rom[19] = 32'b010000000001_01000_101_10111_0010011; // srai x23, x8  -2 >>> 1 = -1
        ///////////////////////////정상작동 여기까지 확인 /////////////////////////////////////


        //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ opcode; // S-Type
        rom[0] = 32'b0000010_00010_00000_000_00010_0100011; // sb x2, 2(x0) [0:7] 32'h0f
        rom[1] = 32'b0000011_00010_00000_001_00011_0100011; // sh x2, 3(x0) [0:15] 32'h4f
        rom[2] = 32'b0000100_00010_00000_010_00100_0100011; // sw x2, 4(x0) [0:31] 32'hff
        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ opcode; // L-Type
        rom[3] = 32'b000000000100_00000_000_00011_0000011; // lb x2, 4(x0); [0:7]
        rom[4] = 32'b000000000100_00000_001_00011_0000011; // lh x3, 4(x0); [0:15]
        rom[5] = 32'b000000000100_00000_010_00011_0000011; // lw x4, 4(x0); [0:31]
        rom[6] = 32'b000000000100_00000_100_00011_0000011; // lbu x5, 4(x0); [0:7] // rdata 분할해야됨 5가지 종류로
        rom[7] = 32'b000000000100_00000_101_00011_0000011; // lhu x6, 4(x0); [0:15]


        //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ opcode; // B-Type 
        rom[0] = 32'b0000000_00010_00010_000_01000_1100011; // beq x2, x2, 8; -> (PC+8) // 참
        rom[1] = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x2, x1 12+11=23 // 미적용
        rom[2] = 32'b0000000_00010_00001_000_01000_1100011; // beq x1, x2, 8; -> (PC+4) // 거짓
        rom[3] = 32'b0100000_00010_00001_000_00100_0110011; // sub x4, x1, x2 11-12=-1 // 적용
        rom[4] = 32'b0000000_00100_00001_001_01000_1100011; // bne x1, x4, 8; -> (PC+8) // 참
        rom[6] = 32'b0000000_00100_00001_100_01000_1100011; // blt x1(11), x4(-1), 8; -> (PC+4) // 거짓
        rom[7] = 32'b0000000_00100_00001_101_01000_1100011; // bge x1(11), x4(-1), 8; -> (PC+imm) // 참
        rom[9] = 32'b0000000_00100_00001_110_01000_1100011; // bltu x1(11), x4(-1), 8; ->  (PC+imm) // 참
        rom[11]= 32'b0000000_00100_00001_111_01000_1100011; // bltu x1(11), x4(-1), 8; ->  (PC+4) // 거짓
        
        //rom[x]=32'b       imm20        _  rd _ opcode; // LU,AU-Type
        rom[0] = 32'b00000000000000000001_00010_0110111; // rd(x2) = 1 << 12 -> 4096
        rom[1] = 32'b00000000000000000001_00010_0010111; // rd(x2) = 4 + 1 << 12 -> 4100
        //rom[x]=32'bimm[20][10:1][11][19:12]_  rd _ opcode; // J-Type
        rom[0] = 32'b0_0000001000_0_00000000__00010_1101111; //  rd = PC + 4, PC += imm -> 4, 16
        rom[4] = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x2, x1
        //rom[x]=32'b imm12      _ rs1 _000_ rd  _ opcode; // JL-Type
        rom[0] = 32'b000000001000_00010_000_00110_1100111; // rd = PC + 4, PC = rs1 + imm -> 4, 24
        rom[6] = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x2, x1
        */
